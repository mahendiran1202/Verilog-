module two_onegatelevel(input i0,i1,s,output y);
 and and_1(a,i0,s);
 and and_2(b.i1,s);
 or or_1(y,a,b);
 endmodule
