




module orgate (a,b,c);
input a,b;
output c;
or or_gate (c,a,b);
endmodule







